module Splice (input [31:0] full_intruc, output [6:0] POC, );


endmodule 